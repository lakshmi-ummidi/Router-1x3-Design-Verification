package router_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	`include "tb_defs.sv"
	`include "source_xtn.sv"
	`include "source_cfg.sv"
	`include "dest_cfg.sv"
	`include "env_cfg.sv"
	`include "s_sequencer.sv"
	`include "s_driver.sv"
	`include "s_monitor.sv"
	`include "source_agt.sv"
	`include "source_agt_top.sv"
	`include "source_seq.sv"
	
	`include "dest_xtn.sv"
	`include "d_sequencer.sv"
	`include "d_driver.sv"
	`include "d_monitor.sv"
	`include "dest_agt.sv"
	`include "dest_agt_top.sv"
	`include "dest_seq.sv"
	
	`include "vsequencer.sv"
	`include "vsequence.sv"
	`include "router_scoreboard.sv"
	`include "env.sv"
	`include "router_test.sv"
	`include "router_vtest.sv"
	
endpackage